library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.game_components.all;
use work.tank_functions.all;
use work.tank_const.all;

entity tank_top_level_tb is
end entity tank_top_level_tb;

architecture testbench of tank_top_level_tb is
	
begin
	
end architecture testbench;