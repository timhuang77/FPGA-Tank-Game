library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.game_components.all;
use work.tank_functions.all;

entity boundary_detection is
	port(
		clk, rst : in std_logic;
		
	);
end entity boundary_detection;

architecture behavioral of boundary_detection is

	
begin
	
	
architecture behavioral;