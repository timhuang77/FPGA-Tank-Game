library IEEE;
use IEEE.std_logic_1164.all;

package tank_const is

	constant TANK_WIDTH : integer := 20;
	constant TANK_HEIGHT : integer := 30;
	constant BULLET_WIDTH : integer := 4;
	constant BULLET_HEIGHT : integer := 8;
	constant TANK_WIDTH_BUFFER : integer := 5;
	
end package tank_const;