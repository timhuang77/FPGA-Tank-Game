library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.game_components.all;
use work.tank_functions.all;

entity game_logic is
	port(
		clk, rst : in std_logic;
		
	);
end entity game_logic;

architecture behavioral of game_logic is

	
begin
	
	
architecture behavioral;